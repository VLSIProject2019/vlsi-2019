// microprocessor